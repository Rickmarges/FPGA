module led_sw(
    output led,
    input sw
);
 
assign led = sw;
 
endmodule